LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;
USE PAKAGEADDER000.ALL;

ENTITY TOPADDER1 IS
	PORT(
		C00, A00, B00 : in std_logic;
		S00, C01 : out std_logic
	);
END TOPADDER1;

ARCHITECTURE TOPADDER01 OF TOPADDER1 IS
SIGNAL SINT1: STD_LOGIC;
SIGNAL CINT1: STD_LOGIC;
SIGNAL CINT2: STD_LOGIC;
BEGIN
	
	US001 : TOPADDER0 PORT MAP(
				A0=>A00,
				B0=>B00,
				S0=>SINT1,
				C0=>CINT1
			);	
		
	US010 : OR0 PORT MAP(
				AI00=>CINT2,
				BI00=>CINT1,
				AO00=>C01
			);
	
	US011 : TOPADDER0 PORT MAP(
				A0=>C00,
				B0=>SINT1,
				S0=>S00,
				C0=>CINT2
			);	
			
END TOPADDER01;