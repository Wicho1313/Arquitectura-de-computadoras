LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;

ENTITY OR0 IS	PORT(
		AI00, BI00 : IN STD_LOGIC;
		AO00 : OUT STD_LOGIC
	);
END OR0;

ARCHITECTURE OR00 OF OR0 IS 
	BEGIN
		AO00<=AI00 OR BI00;
	END ARCHITECTURE;
		