LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;

PACKAGE PACKAGEMUL00 IS
	COMPONENT AND0
		PORT(
			AI00, BI00 : IN STD_LOGIC;
			AO00 : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT TOPADDER1
		PORT(
			C00, A00, B00 : in std_logic;
			S00, C01 : out std_logic
		);
	END COMPONENT;
END PACKAGEMUL00;