LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;

PACKAGE PAKAGEADDER000 IS
	COMPONENT TOPADDER0 
		PORT(
			A0, B0 : in std_logic;
			S0, C0 : out std_logic
		);
	END COMPONENT;
	
	COMPONENT OR0
		PORT(
			AI00, BI00 : IN STD_LOGIC;
			AO00 : OUT STD_LOGIC
		);
	END COMPONENT;
END PAKAGEADDER000;