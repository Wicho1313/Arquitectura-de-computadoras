LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;

PACKAGE pakaguecom00 IS
	COMPONENT AND0
		PORT(
			AI00, BI00 : IN STD_LOGIC;
			AO00 : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT OR0
		PORT(
			AI00, BI00 : IN STD_LOGIC;
			AO00 : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT NOT0
		PORT(
			AI00 : IN STD_LOGIC;
			AO00 : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT XOR0
		PORT(
			AI00, BI00 : IN STD_LOGIC;
			AO00 : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT NAND0
		PORT(
			AI00, BI00 : IN STD_LOGIC;
			AO00 : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT NOR0
		PORT(
			AI00, BI00 : IN STD_LOGIC;
			AO00 : OUT STD_LOGIC
		);
	END COMPONENT;
	
	COMPONENT XNOR0
		PORT(
			AI00, BI00 : IN STD_LOGIC;
			AO00 : OUT STD_LOGIC
		);
	END COMPONENT;
	
END pakaguecom00;